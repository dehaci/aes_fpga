----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 2018/05/09 18:36:19
-- Design Name: 
-- Module Name: keyexpansion - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity keyexpansion is
	port(
			clk : in std_logic;
			original_key : in std_logic_vector(0 to 127);

			round0 : out std_logic_vector(0 to 127);
			round1 : out std_logic_vector(0 to 127);
			round2 : out std_logic_vector(0 to 127);
			round3 : out std_logic_vector(0 to 127);
			round4 : out std_logic_vector(0 to 127);
			round5 : out std_logic_vector(0 to 127);
			round6 : out std_logic_vector(0 to 127);
			round7 : out std_logic_vector(0 to 127);
			round8 : out std_logic_vector(0 to 127);
			round9 : out std_logic_vector(0 to 127);
			round10 : out std_logic_vector(0 to 127)
		);
end keyexpansion;

architecture Behavioral of keyexpansion is
	type array_2d is array (0 to 15, 0 to 15) of std_logic_vector(7 downto 0);
	type array_1d is array (1 to 10) of std_logic_vector(31 downto 0);
	constant lut : array_2d :=
	(
	  ---- 0 ---- 1 ---- 2 ---- 3 ---- 4 ---- 5 ---- 6 ---- 7 ---- 8 ---- 9 ---- A ---- B ---- C ---- D ---- E ---- F ----
    	(x"63", x"7C", x"77", x"7B", x"F2", x"6B", x"6F", x"C5", x"30", x"01", x"67", x"2B", x"FE", x"D7", x"AB", x"76"),  -- 0 --
		(x"CA", x"82", x"C9", x"7D", x"FA", x"59", x"47", x"F0", x"AD", x"D4", x"A2", x"AF", x"9C", x"A4", x"72", x"C0"),  -- 1 --      
		(x"B7", x"FD", x"93", x"26", x"36", x"3F", x"F7", x"CC", x"34", x"A5", x"E5", x"F1", x"71", x"D8", x"31", x"15"),  -- 2 --
		(x"04", x"C7", x"23", x"C3", x"18", x"96", x"05", x"9A", x"07", x"12", x"80", x"E2", x"EB", x"27", x"B2", x"75"),  -- 3 --
		(x"09", x"83", x"2C", x"1A", x"1B", x"6E", x"5A", x"A0", x"52", x"3B", x"D6", x"B3", x"29", x"E3", x"2F", x"84"),  -- 4 --
		(x"53", x"D1", x"00", x"ED", x"20", x"FC", x"B1", x"5B", x"6A", x"CB", x"BE", x"39", x"4A", x"4C", x"58", x"CF"),  -- 5 --
		(x"D0", x"EF", x"AA", x"FB", x"43", x"4D", x"33", x"85", x"45", x"F9", x"02", x"7F", x"50", x"3C", x"9F", x"A8"),  -- 6 --
		(x"51", x"A3", x"40", x"8F", x"92", x"9D", x"38", x"F5", x"BC", x"B6", x"DA", x"21", x"10", x"FF", x"F3", x"D2"),  -- 7 --
		(x"CD", x"0C", x"13", x"EC", x"5F", x"97", x"44", x"17", x"C4", x"A7", x"7E", x"3D", x"64", x"5D", x"19", x"73"),  -- 8 --
		(x"60", x"81", x"4F", x"DC", x"22", x"2A", x"90", x"88", x"46", x"EE", x"B8", x"14", x"DE", x"5E", x"0B", x"DB"),  -- 9 --
		(x"E0", x"32", x"3A", x"0A", x"49", x"06", x"24", x"5C", x"C2", x"D3", x"AC", x"62", x"91", x"95", x"E4", x"79"),  -- A --
		(x"E7", x"C8", x"37", x"6D", x"8D", x"D5", x"4E", x"A9", x"6C", x"56", x"F4", x"EA", x"65", x"7A", x"AE", x"08"),  -- B --
		(x"BA", x"78", x"25", x"2E", x"1C", x"A6", x"B4", x"C6", x"E8", x"DD", x"74", x"1F", x"4B", x"BD", x"8B", x"8A"),  -- C --
		(x"70", x"3E", x"B5", x"66", x"48", x"03", x"F6", x"0E", x"61", x"35", x"57", x"B9", x"86", x"C1", x"1D", x"9E"),  -- D --
		(x"E1", x"F8", x"98", x"11", x"69", x"D9", x"8E", x"94", x"9B", x"1E", x"87", x"E9", x"CE", x"55", x"28", x"DF"),  -- E --
		(x"8C", x"A1", x"89", x"0D", x"BF", x"E6", x"42", x"68", x"41", x"99", x"2D", x"0F", x"B0", x"54", x"BB", x"16")   -- F --
	);
	constant rcon : array_1d :=
	(
		x"01000000",
		x"02000000",
		x"04000000",
		x"08000000",
		x"10000000",
		x"20000000",
		x"40000000",
		x"80000000",
		x"1b000000",
		x"36000000"
	);
begin
	process(clk)
		variable all_w : std_logic_vector(0 to 1407) := (others => '0');
		variable temp : std_logic_vector(0 to 31) := (others => '0');
		variable temp1 : std_logic_vector(0 to 31) := (others => '0');
		variable temp2 : std_logic_vector(0 to 31) := (others => '0');
		variable temp3 : std_logic_vector(0 to 31) := (others => '0');
		begin
			if rising_edge(clk) then
				all_w(0 to 127) := original_key;
					for i in 4 to 43 loop
						temp := all_w((i-1)*32 to (i-1)*32+31);
						if i-(i/4)*4 = 0 then
							temp1 := temp(8 to 31) & temp(0 to 7);
							for n in 0 to 3 loop
								temp2(n*8 to n*8+7) := lut(conv_integer(temp1(n*8 to n*8+3)),conv_integer(temp1(n*8+4 to n*8+7)));
							end loop;
							temp3 := temp2 xor rcon(i/4);
							all_w(i*32 to i*32+31) := temp3 xor all_w((i-4)*32 to (i-4)*32+31);
						else
							all_w(i*32 to i*32+31) := temp xor all_w((i-4)*32 to (i-4)*32+31);
						end if;
					end loop;
					round0 <= all_w(0 to 127);
					round1 <= all_w(128 to 255);
					round2 <= all_w(256 to 383);
					round3 <= all_w(384 to 511);
					round4 <= all_w(512 to 639);
					round5 <= all_w(640 to 767);
					round6 <= all_w(768 to 895);
					round7 <= all_w(896 to 1023);
					round8 <= all_w(1024 to 1151);
					round9 <= all_w(1152 to 1279);
					round10 <= all_w(1280 to 1407);
			end if;
	end process;

end Behavioral;
